module top
(
);