module IDE

(
input [31:0] instruction;
outpu 